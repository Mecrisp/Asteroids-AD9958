
`default_nettype none

/* verilator lint_off UNUSEDSIGNAL */

module fiftyfivenm_rublock(
    input wire rconfig,
    input wire clk,
    input wire rsttimer,
    input wire shiftnld,
    input wire captnupdt,
    input wire regin,
    output wire regout
  );

  assign regout = 0;



endmodule

/* verilator lint_on UNUSEDSIGNAL */
